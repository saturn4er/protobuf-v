module wiretest
